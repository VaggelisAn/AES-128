/**         Implementation of the AES-128 Encryptor     **/
/**                 Key Expansion Module                **/
/** Vaggelis Ananiadis 03409, Nikh-Maria Kalantzh 03502 **/

/*
Key Expansion Algorithm explanation:
From: https://engineering.purdue.edu/kak/compsec/NewLectures/Lecture8.pdf

Let the four words of the round key for the ith round be:
wi, wi+1, wi+2, wi+3
for example round1 (i=1*4) : w4, w5, w6, w7,
round2 (i=2*4) : w8, w9, w10, w11 etc.  

We have:
wi+5 = wi+4 (+) wi+1
wi+6 = wi+5 (+) wi+2
wi+7 = wi+6 (+) wi+3

Now we need to figure out wi+4, obtained by:
wi+4 = wi (+) g(wi+3),

g(w) consists of the following steps: (w is a word)
1. One byte left circular rotation of w
2. Byte substitution for each of the four bytes of w, using the sbox table from SubBytes
3. XOR the obtained bytes with the round constant for the ith round, Rcon[i].

Τhe Round Constant, Rcon, is a word whose three rightmost bytes are always zero
Rcon[i] = [RC[i], 0x00, 0x00, 0x00], where RC[i] is calculated through a recursion, as follows:
RC[1] = 0x01
RC[j] = 0x02 * RC[j-1]
This steps destroys any symmetries that may have been introduced in other steps in the key expansion algo
*/

`timescale 1ns / 1ps
//`include "lut//sbox.v" is not used due to coding problems explained below

module KeyExpansion(key, RoundKeys);
input [127:0] key;
output reg [1407:0] RoundKeys;

reg [31:0] w [0:43];

reg [31:0] rot;
reg [31:0] subword;
reg [31:0] rcon;

integer i;

`include "sbox.v"

always@* begin
    w[0] = key[127:96];
    w[1] = key[95:64];
    w[2] = key[63:32];
    w[3] = key[31:0];
    #5;
    for (i = 4; i < 44; i = i + 1) begin : keyExpLoop
        if (i % 4 == 0) begin
            rot = rot_w(w[i - 1]);
            subword[31:24] = sbox(rot[31:24]);
            subword[23:16] = sbox(rot[23:16]);
            subword[15:8] = sbox(rot[15:8]);
            subword[7:0] = sbox(rot[7:0]);
            rcon = rcon_w(i>>2); // divide by 4
            w[i] = w[i - 4] ^ subword ^ rcon;

            //$display("w[i - 1]=%h", w[i - 1]);
            //$display("subword=%h", subword);
            //$display("rcon=%h", rcon);
            //$display("w[%h]=%h",i, w[i]);
        end 
        else
            w[i] = w[i - 4] ^ w[i - 1];
            //$display("w[%h]=%h",i, w[i]);
    #5; // simulate delay so we can monitor results in gtkwave
    end

    RoundKeys = {w[0], w[1], w[2], w[3], w[4], w[5], w[6], w[7],
                w[8], w[9], w[10], w[11], w[12], w[13], w[14], w[15],
                w[16], w[17], w[18], w[19], w[20], w[21], w[22], w[23],
                w[24], w[25], w[26], w[27], w[28], w[29], w[30], w[31],
                w[32], w[33], w[34], w[35], w[36], w[37], w[38], w[39],
                w[40], w[41], w[42], w[43]};

end

function [31:0] rot_w;
    input [31:0] word;
    rot_w = {word[23:0], word[31:24]};;
endfunction

// As generated by our generate_rcon.py script:
function [31:0] rcon_w;
	input[3:0] round;
    begin
    case(round)	
        4'h1: rcon_w=32'h01000000;
        4'h2: rcon_w=32'h02000000;
        4'h3: rcon_w=32'h04000000;
        4'h4: rcon_w=32'h08000000;
        4'h5: rcon_w=32'h10000000;
        4'h6: rcon_w=32'h20000000;
        4'h7: rcon_w=32'h40000000;
        4'h8: rcon_w=32'h80000000;
        4'h9: rcon_w=32'h1b000000;
        4'hA: rcon_w=32'h36000000;
        default: rcon_w=32'h00000000;
    endcase
    end 
endfunction	

endmodule